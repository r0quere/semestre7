
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.all;

--/////////////////////
--    A COMPLETER
--/////////////////////